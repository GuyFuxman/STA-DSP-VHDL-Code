-- FFT.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity FFT is
	port (
		fft_ii_0_clk_clk              : in  std_logic                     := '0';             --    fft_ii_0_clk.clk
		fft_ii_0_rst_reset_n          : in  std_logic                     := '0';             --    fft_ii_0_rst.reset_n
		fft_ii_0_sink_valid           : in  std_logic                     := '0';             --   fft_ii_0_sink.valid
		fft_ii_0_sink_ready           : out std_logic;                                        --                .ready
		fft_ii_0_sink_error           : in  std_logic_vector(1 downto 0)  := (others => '0'); --                .error
		fft_ii_0_sink_startofpacket   : in  std_logic                     := '0';             --                .startofpacket
		fft_ii_0_sink_endofpacket     : in  std_logic                     := '0';             --                .endofpacket
		fft_ii_0_sink_data            : in  std_logic_vector(47 downto 0) := (others => '0'); --                .data
		fft_ii_0_source_valid         : out std_logic;                                        -- fft_ii_0_source.valid
		fft_ii_0_source_ready         : in  std_logic                     := '0';             --                .ready
		fft_ii_0_source_error         : out std_logic_vector(1 downto 0);                     --                .error
		fft_ii_0_source_startofpacket : out std_logic;                                        --                .startofpacket
		fft_ii_0_source_endofpacket   : out std_logic;                                        --                .endofpacket
		fft_ii_0_source_data          : out std_logic_vector(46 downto 0)                     --                .data
	);
end entity FFT;

architecture rtl of FFT is
	component FFT_fft_0 is
		port (
			clk          : in  std_logic                     := 'X';             -- clk
			reset_n      : in  std_logic                     := 'X';             -- reset_n
			sink_valid   : in  std_logic                     := 'X';             -- valid
			sink_ready   : out std_logic;                                        -- ready
			sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			sink_sop     : in  std_logic                     := 'X';             -- startofpacket
			sink_eop     : in  std_logic                     := 'X';             -- endofpacket
			inverse      : in  std_logic                     := 'X';             -- data
			fftpts_in    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- data
			sink_imag    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			sink_real    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			source_valid : out std_logic;                                        -- valid
			source_ready : in  std_logic                     := 'X';             -- ready
			source_error : out std_logic_vector(1 downto 0);                     -- error
			source_sop   : out std_logic;                                        -- startofpacket
			source_eop   : out std_logic;                                        -- endofpacket
			fftpts_out   : out std_logic_vector(14 downto 0);                    -- data
			source_imag  : out std_logic_vector(15 downto 0);                    -- data
			source_real  : out std_logic_vector(15 downto 0)                     -- data
		);
	end component FFT_fft_0;

	signal fft_0_source_imag : std_logic_vector(15 downto 0); -- port fragment
	signal fft_0_source_real : std_logic_vector(15 downto 0); -- port fragment
	signal fft_0_fftpts_out  : std_logic_vector(14 downto 0); -- port fragment

begin

	fft_0 : component FFT_fft_0
		port map (
			clk                      => fft_ii_0_clk_clk,                 --    clk.clk
			reset_n                  => fft_ii_0_rst_reset_n,             --    rst.reset_n
			sink_valid               => fft_ii_0_sink_valid,              --   sink.valid
			sink_ready               => fft_ii_0_sink_ready,              --       .ready
			sink_error               => fft_ii_0_sink_error,              --       .error
			sink_sop                 => fft_ii_0_sink_startofpacket,      --       .startofpacket
			sink_eop                 => fft_ii_0_sink_endofpacket,        --       .endofpacket
			sink_real(15 downto 0)   => fft_ii_0_sink_data(47 downto 32), --       .data
			sink_imag(15 downto 0)   => fft_ii_0_sink_data(31 downto 16), --       .data
			fftpts_in(14 downto 0)   => fft_ii_0_sink_data(15 downto 1),  --       .data
			inverse                  => fft_ii_0_sink_data(0),            --       .data
			source_valid             => fft_ii_0_source_valid,            -- source.valid
			source_ready             => fft_ii_0_source_ready,            --       .ready
			source_error             => fft_ii_0_source_error,            --       .error
			source_sop               => fft_ii_0_source_startofpacket,    --       .startofpacket
			source_eop               => fft_ii_0_source_endofpacket,      --       .endofpacket
			source_real(15 downto 0) => fft_0_source_real(15 downto 0),   --       .data
			source_imag(15 downto 0) => fft_0_source_imag(15 downto 0),   --       .data
			fftpts_out(14 downto 0)  => fft_0_fftpts_out(14 downto 0)     --       .data
		);

	fft_ii_0_source_data <= fft_0_source_real(15 downto 0) & fft_0_source_imag(15 downto 0) & fft_0_fftpts_out(14 downto 0);

end architecture rtl; -- of FFT
