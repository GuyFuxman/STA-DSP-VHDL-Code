/* 
RON KRAKOVSKY
Convolution with hann function, window function.
*/

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--------------------------------------------------

entity Window_Multipication is
generic(
	samples : integer := 512;
	width_input_data_bits : integer := 10; 
	width_memory_data : integer := 10 -- ufix10_En8
);
port(	
	csi_sink_clk	 	 : in std_logic; -- clock
	rsi_sink_reset	 	 : in std_logic; -- reset in LOW = '0'
	asi_sink_valid_data	 : in std_logic; -- valid for start convolution, start when fft need for data.(start of pucket)
	asi_sink_data		 : in std_logic_vector(width_input_data_bits - 1 downto 0); -- s10_En0 ,input data 
	aso_source_data		 : out std_logic_vector(width_input_data_bits - 1 downto 0); -- s10_En0 ,output data
	aso_Window_Multipication : out std_logic

);
end Window_Multipication;  

--------------------------------------------------

architecture arch_Window_Multipication of Window_Multipication is
type mem_t is array(0 to samples-1) of unsigned(width_memory_data-1 downto 0); -- ufix10_En8
signal ram : mem_t;
attribute ram_init_file : string;
attribute ram_init_file of ram :
signal is "Hann1024.mif";

TYPE STATE_TYPE IS (idle, start);
signal state : STATE_TYPE;

signal s_convolution : integer;
signal index_hann : integer range 0 to samples;
begin

    process(csi_sink_clk, rsi_sink_reset)
    begin
		if rsi_sink_reset = '0' then 
			s_convolution <= 0;
			index_hann <= 0;
			state <= idle;
			aso_Window_Multipication <= '0';
		elsif rising_edge(csi_sink_clk) then 
			case state is 
				when idle => 
					s_convolution <= 0;
					index_hann <= 0;
					if asi_sink_valid_data = '1' then
						state <= start;
						aso_Window_Multipication <= '1';
					end if;
					
				when start => 
					if index_hann = samples - 2 then 
						index_hann <= 0;
						state <= idle;
					else
						s_convolution <= to_integer(ram(index_hann)) * to_integer(signed(asi_sink_data));
						index_hann <= index_hann + 1;
						if asi_sink_valid_data = '1' then
							index_hann <= 0;
						end if;
						
					end if;
			end case;	
		end if;
    end process;
aso_source_data <= std_logic_vector(to_signed(s_convolution/256,width_input_data_bits)); -- 2^8 because we dont need fix point number
end arch_Window_Multipication;
